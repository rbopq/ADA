----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    22:43:23 05/07/2016 
-- Design Name: 
-- Module Name:    multiplicador_mux-2_1 - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity multiplicador_mux_2_1 is
	Port(operando_1 : in STD_LOGIC_VECTOR(0 downto 0);
		 operando_2 : in STD_LOGIC_VECTOR(0 downto 0);
		 sel        : in STD_LOGIC_VECTOR(0 downto 0));
end multiplicador_mux_2_1;

architecture Behavioral of multiplicador_mux_2_1 is
begin
end Behavioral;

